module siso (
    clk,clear,si,so
);
    input clk,clear,si;
    output so;
    reg [3:0]tmp;
    
    
endmodule